--###############################
--# Project Name : 
--# File         : 
--# Project      : VHDL RAM model
--# Engineer     : 
--# Modification History
--###############################
-- VHDL model for altera

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;

ENTITY dp16x16 IS
	PORT
	(
		address_a	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		address_b	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		clock_a		: IN STD_LOGIC  := '1';
		clock_b		: IN STD_LOGIC 	:= '1';
		data_a		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data_b		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		wren_a		: IN STD_LOGIC  := '0';
		wren_b		: IN STD_LOGIC  := '0';
		q_a			: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		q_b			: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END dp16x16;

architecture rtl of dp16x16 is
	constant ram_depth : natural := 16;
	constant ram_width : natural := 16;
	type memory is array(0 to ram_depth-1) of std_logic_vector(ram_width-1 downto 0);
	impure function init_mem return memory is
		file afile : text open read_mode is "dp16x16.dat";
		variable aline : line;
		variable amem : memory;
		variable bv : bit_vector(ram_width-1 downto 0);
	begin
		for i in 0 to ram_depth-1 loop
			readline(afile,aline);
			read(aline,bv);
			amem(i) := To_StdLogicVector(bv);
		end loop;
		return amem;
	end function;
	shared variable mem : memory := init_mem;
begin
	RAM_A : process(clock_a)
	begin
		if (clock_a'event and clock_a='1') then
				if (wren_a = '0') then
					q_a <= mem(to_integer(unsigned(address_a)));
				else
					mem(to_integer(unsigned(address_a))) := data_a;
					q_a <= data_a;  -- ????
				end if;
		end if;
	end process RAM_A;
	
	RAM_B : process(clock_b)
	begin
		if (clock_b'event and clock_b='1') then
				if (wren_b = '0') then
					q_b <= mem(to_integer(unsigned(address_b)));
				else
					mem(to_integer(unsigned(address_b))) := data_b;
					q_b <= data_b;  -- ????
				end if;
		end if;
	end process RAM_B;
	
	
end rtl;
